magic
tech sky130A
magscale 1 2
timestamp 1713442895
<< metal1 >>
rect 104 1610 304 1810
rect 114 802 314 1002
use sky130_fd_pr__res_generic_po_4WEV9M  R1
timestamp 1713442895
transform 1 0 213 0 1 1308
box -266 -761 266 761
<< labels >>
flabel metal1 114 802 314 1002 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 104 1610 304 1810 0 FreeSans 256 0 0 0 VSS
port 1 nsew
<< end >>
