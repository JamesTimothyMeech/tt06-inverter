** sch_path: /home/james/Desktop/TinyTapeout/TinyTapeoutAnalog/tt06-inverter/xschem/inverter.sch
.subckt inverter VDD VSS
*.PININFO VDD:B VSS:B
XR1 VSS VDD VSS sky130_fd_pr__res_high_po_0p35 L=0.35 mult=1 m=1
.ends
.end
