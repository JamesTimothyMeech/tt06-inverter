** sch_path: /home/james/Desktop/TinyTapeout/TinyTapeoutAnalog/tt06-inverter/xschem/inverter.sch
.subckt inverter VDD VSS
*.PININFO VDD:B VSS:B
R1 VSS VDD sky130_fd_pr__res_generic_po W=1 L=1 m=1
.ends
.end
